library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;


entity i2s_delay_line is
port (
    clk : std_logic;
    reset : std_logic 
);
end entity;

architecture rtl of i2s_delay_line is
begin

end architecture;

